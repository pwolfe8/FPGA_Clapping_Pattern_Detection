--Engineer     : Philip Wolfe
--Date         : 11/30/2017
--Name of file : Top_Level_Detector.vhd
--Description  : Top level clapping pattern detector file.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Top_Level_Detector is
    port (
        -- inputs --
        _name_		: in  _type_;
        -- outputs --
        _name_		: out _type_
    );
end Top_Level_Detector;

architecture Top_Level_Detector_arch of Top_Level_Detector is
    -- constant definitions
    
    -- signal declarations
    

begin
    
    
end Top_Level_Detector_arch;
