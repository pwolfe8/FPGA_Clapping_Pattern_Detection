will@Kira.30855:1511711835